module planner

