module main
// const version = '1.0.21'

//TODO: NOT WORKING,WHY?
