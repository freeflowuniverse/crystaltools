module builder

