module libp2p


// println(redis.get("test"))

