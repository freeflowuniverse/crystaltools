module ct

pub const version = '1.0.21'

