module manifestor
import os

struct ExecutorLocal{
}


