module tfgrid


struct Tags {
	tags Tag[]
}

struct Tag {
	key string
	val string
}


