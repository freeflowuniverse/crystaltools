module installerpublisher
