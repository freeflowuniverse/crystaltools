module manifestor
import os


