	
	
module main
// import despiegk.crystallib.
import os

fn main() {


}