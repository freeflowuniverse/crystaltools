	
	
module main
import despiegk.crystallib.imagemagick
import os


fn main() {
	mut magic := imagemagick.new()
	magic.add("") or {panic("did not load")}
	// println(magic)

	magic.downsize("/Users/despiegk/code/github/threefoldfoundation/info_threefold_pub/wiki/","/Users/despiegk/backup_images/threefold/") or {panic("could not downsize. $err")}


	
	
}