module config
// import gittools

pub struct ConfigData {
pub mut:
}

