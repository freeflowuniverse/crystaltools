	
	
module main
// import freeflowuniverse.crystallib.
import os

fn main() {


}