module docker

//build ssh enabled alpine docker image
//has default ssh key in there
// pub fn (mut e DockerEngine) builder_build() ?DockerImage {

// 	//TODO: create temporary directory
// 	// store the docker file & the boot.sh file
// 	// run the docker builder
// 	// return the image which has been build

// 	//use template engine to get the base in
// 	base = "alpine:3.13"
// 	redis_enable = false

// 	//template engine/write files ... (use variables)


// }


//if docker image for builder not build yet (locally, then do so) 
//start a container with the image of the builder
//do a test that ssh is working with predefined key
// pub fn (mut e DockerEngine) builder_container_get(name:string) ?DockerContainer {


// }

