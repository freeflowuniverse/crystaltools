module tmux

import os
import vredis2
import builder

struct Tmux {
mut:
	sessions map[string]Session
	node     builder.Node
}

pub fn new(args builder.NodeArguments) Tmux {
	mut t := Tmux{
		sessions: map[string]Session{}
		node: builder.node_get(args) or { panic(err) }
	}
	os.log('scan')
	t.scan()
	return t
}

pub fn (mut t Tmux) session_get(name string, restart bool) Session {
	name_l := name.to_lower()
	mut session := Session{}
	if name_l in t.sessions {
		session = t.sessions[name_l]
	} else {
		session = init_session(t, name_l)
		t.sessions[name_l] = session
	}
	if restart {
		session.restart()
	}
	return session
}

pub fn (mut t Tmux) scan() {
	exec_list := t.node.executor.exec('tmux list-sessions') or { '1' }

	if exec_list == '1' {
		// No server running
		return
	}

	mut done := map[string]bool{}

	out := t.node.executor.exec("tmux list-windows -a -F '#{session_name}|#{window_name}|#{window_id}|#{pane_active}|#{pane_pid}|#{pane_start_command}'") or {
		panic("Can't execute")
	}
	for line in out.split_into_lines() {
		if line.contains('|') {
			line_arr := line.split('|')
			session_name := line_arr[0]
			window_name := line_arr[1]
			window_id := line_arr[2]
			pane_active := line_arr[3]
			pane_pid := line_arr[4]
			pane_start_command := line_arr[5] or { '' }

			key := session_name + '-' + window_name
			os.log(' - found session: $session_name $window_name id: $window_id $pane_active, $pane_pid, $pane_start_command')
			mut session := t.session_get(session_name, false)
			window_name_l := window_name.to_lower()

			if key in done {
				error('Duplicated window name: $key')
			}
			mut active := false
			if pane_active == '1' {
				active = true
			}
			if window_name != 'notused' {
				mut window := session.window_get(window_name_l)
				window.id = (window_id.replace('@', '')).int()
				window.pid = pane_pid.int()
				window.active = active
				done[key] = true
			}
			t.sessions[session_name] = session
		}
	}
}

pub fn (mut t Tmux) stop() {
	for _, mut session in t.sessions {
		session.stop()
	}
	mut redis := vredis2.connect('localhost:6379') or { panic("Couldn't connect to redis client") }
	redis.del('tmux:active_session') or { 1 }
	redis.del('tmux:active_window') or { 1 }
}

pub fn (mut t Tmux) list() {
	for _, session in t.sessions {
		for _, window in session.windows {
			println('- $session.name: $window.name')
		}
	}
}
