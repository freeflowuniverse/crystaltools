module publishingtools

import os

// nothing kept in mem, just to process one iteration
struct PageActor {
pub mut:
	page      Page
	page_errors map[string][]PageError // page_errors[page.path]
	site      Site
	publtools PublTools
}

// return fullpath,pageobject
pub fn (site Site) pageactor_get(name string, publtools PublTools) ?PageActor {
	namelower := name_fix(name)
	if namelower in site.pages {
		page := site.pages[namelower]
		return PageActor{
			page: page // {page|errors:page.errors.clone()}
			publtools: publtools
			site: site
		}
	}
	return error('Could not find page $namelower in site $site.name')
}

pub fn (pageactor PageActor) path_get() string {
	return os.join_path(pageactor.site.path, pageactor.page.path)
}

// will load the content, check everything, return true if ok
pub fn (mut pageactor PageActor) check() bool {
	//content := pageactor.markdown_get()
	if pageactor.page.state == PageStatus.error {
		return false
	}
	return true
}

// process the markdown content and include other files, find links, ...
// the content is the processed 
// originSite is the site that wants to include a markdown page
pub fn (mut pageactor PageActor) markdown_get(originSite string) string {
	if pageactor.page.content != '' {
		// means was already processed, if fast enough we can leave this away that way we know includes are dynamic
		return pageactor.page.content
	}
	mut content := pageactor.markdown_load() or { panic(err) }
	// for i in 0 .. 10 {
	// 	if i>9 {
	// 		panic ("too many level of includes in ${pageactor.path_get()}")
	// 	}
	// 	if i>3{
	// 		panic("seems off, need to first find why the uncludes don't get replaced")
	// 	}		
	content = pageactor.process_includes(content) // should be recursive now
	// 	if !content.contains("!!!include") {
	// 		//means we got all the includes 
	// 		break
	// 	}
	// 	// println( content)
	// }
	//if pageactor.page.errors.len > 0 {
	if pageactor.page_errors[pageactor.page.path].len > 0 {
		pageactor.page.state = .error
	}
	// check for links
	mut res := link_parser(content)
	// mut link:=Link{}
	for mut link in res.links {
		content = link.check_replace(content, mut pageactor.publtools, mut pageactor.site, originSite)
		// println("${replaceaction.original_text}->${replaceaction.new_text}")
		if link.state == LinkState.notfound {
			mut cat := PageErrorCat.brokenlink
			if link.cat == LinkType.image {
				cat = PageErrorCat.brokenimage
			}
			page_error := PageError{
				line: ''
				linenr: 0
				msg: link.error_msg_get()
				cat: cat
			}
			pageactor.error_add(page_error)
		}
	}
	pageactor.page.content = content
	return pageactor.page.content
}

pub fn (pageactor PageActor) markdown_load() ?string {
	// path_surce2 := pageactor.path_get()
	content := os.read_file(pageactor.path_get()) or {
		path_source := pageactor.path_get()
		println('Failed to open $path_source')
		return err
	}
	return content
}

pub fn (mut pageactor PageActor) error_add(error PageError) {
	if pageactor.page.state != PageStatus.error {
		// only add when not in error mode yet, because means check was already done
		//pageactor.page.errors << error
		pageactor.page_errors[pageactor.page.path] << error
	}
	println(' ** ERROR: in file $pageactor.path_get()')
	println(error)
}

fn (mut pageactor PageActor) process_includes(content string) string {
	mut lines := ''
	mut nr := 0
	for line in content.split_into_lines() {
		// println (line)
		nr++
		mut linestrip := line.trim(' ')
		if linestrip.starts_with('!!!include') {
			name := linestrip['!!!include'.len + 1..]
			mut pt := pageactor.publtools
			mut pageactor_linked := pt.page_get(name) or {
				page_error := PageError{
					line: line
					linenr: nr
					msg: "Cannot inlude '$name'\n$err"
					cat: PageErrorCat.brokeninclude
				}
				pageactor.error_add(page_error)
				lines += '> ERROR: $page_error.msg'
				continue
			}
			if pageactor_linked.path_get() == pageactor.path_get() {
				panic('recursive include: $pageactor_linked.path_get()')
			}
			pageactor_linked.page.nrtimes_inluded++
			// path11 := pageactor_linked.page
			content_linked := pageactor_linked.markdown_get(pageactor.site.name)
			lines += content_linked + '\n'
		} else {
			lines += line + '\n'
		}
	}
	return lines
}
